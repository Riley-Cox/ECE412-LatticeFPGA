// Defines for Upduino
//`define SPI_FLASH
`define INTERNAL_OSC
